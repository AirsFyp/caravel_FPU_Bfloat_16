module FPU_dec_ctl (
input fpu_active,
input [31:0] instr,
output [114:0] out 
);

wire [31:0] i;
assign i[31:0] = (fpu_active) ? instr[31:0] : {32{1'b0}};

localparam rs1 	= 0;
localparam rs2 	= 1;
localparam rd  	= 2;
localparam vs1 	= 3;
localparam vs2 	= 4;
localparam vs3 	= 5;
localparam vd  	= 6;
localparam imm12 	= 7;
localparam simm  	= 8;
localparam vm    	= 9;
localparam vsetvl 	= 10;
localparam valu   	= 11;
localparam vmul   	= 12;
localparam vdiv   	= 13;
localparam vrem   	= 14;
localparam vlsu   	= 15;
localparam vload  	= 16;
localparam vstore 	= 17;
localparam vadd   	= 18;
localparam vsub   	= 19;
localparam vand   	= 20;
localparam vor    	= 21;
localparam vxor   	= 22;
localparam vsll   	= 23;
localparam vsra   	= 24;
localparam vsrl   	= 25;
localparam vmslt  	= 26;
localparam vmseq  	= 27;
localparam vmsne  	= 28;
localparam vmsle  	= 29;
localparam vmsgt  	= 30;
localparam unsign   	= 31;
localparam sign  	= 32;
localparam by  	= 33;
localparam half         = 34;
localparam word         = 35;
localparam element      = 36;
localparam csr_read     = 37;
localparam csr_write_1  = 38;
localparam csr_write_2  = 39;
localparam rs1_sign     = 40;
localparam rs2_sign     = 41;
localparam vs1_sign     = 42;
localparam vs2_sign     = 43;
localparam low          = 44;
localparam unit_st      = 45;
localparam stride       = 46;
localparam indexed      = 47;
localparam zero_extend  = 48;
localparam sign_extend  = 49;
localparam i0_only      = 50;
localparam legal        = 51;
localparam vmin         = 52;
localparam vmax         = 53;
localparam fs1          = 54;
localparam fs2          = 55;
localparam fs3          = 56;
localparam fd           = 57;
localparam vfadd        = 58;
localparam vfsub        = 59;
localparam vfmin        = 60;
localparam vfmax        = 61;
localparam vfmv         = 62;
localparam vmfeq        = 63;
localparam vmfle        = 64;
localparam vmflt        = 65;
localparam vmfne        = 66;
localparam vmfgt        = 67;
localparam vmfge        = 68;
localparam vfdiv        = 69;
localparam vfmul        = 70;
localparam vfmadd       = 71;
localparam vfmsub       = 72;
localparam vfsqrt       = 73;
localparam vfpu         = 74;
localparam fadd         = 75;
localparam fsub         = 76;
localparam fmul         = 77;
localparam fdiv         = 78;
localparam fsqrt        = 79;
localparam fmin         = 80;
localparam fmax         = 81;
localparam fmvx         = 82;
localparam fmvf         = 83;
localparam feq          = 84;
localparam flt          = 85;
localparam fle          = 86;
localparam fmadd        = 87;
localparam fmsub        = 88;
localparam single_p     = 89;
localparam double_p     = 90;
localparam half_p       = 91;
localparam scalar_fpu   = 92;
localparam vector_fpu   = 93;
localparam vfmvs        = 94;
localparam vfmvf        = 95;
localparam vfcvt_x_f    = 96;
localparam vfcvt_f_x    = 97;
localparam fcvt_w_p     = 98;
localparam fcvt_p_w     = 99;
localparam fnmsub       = 100;
localparam fnmadd       = 101;
localparam fsgnj        = 102;
localparam fsgnjn       = 103;
localparam fsgnjx       = 104;
localparam fclass       = 105;
localparam vfnmadd      = 106;
localparam vfnmsub      = 107;
localparam vfsgnj       = 108;
localparam vfsgnjn      = 109;
localparam vfsgnjx      = 110;
localparam vfclass      = 111;
localparam flsu         = 112;
localparam fload        = 113;
localparam fstore       = 114;

assign out[rs1] = (!i[30]&!i[29]&i[28]&!i[27]&i[26]&i[25]&i[14]&!i[13]&!i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[29]&!i[28]&i[27]&i[25]
    &i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]
    &i[29]&!i[28]&i[26]&i[25]&i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (i[31]&i[30]&i[28]&!i[27]&!i[25]&!i[24]&!i[23]
    &!i[22]&!i[21]&!i[20]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]
    &i[1]&i[0]) | (i[31]&i[30]&i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]
    &!i[21]&!i[20]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]
    &i[0]) | (i[31]&i[30]&!i[29]&i[28]&!i[27]&!i[25]&!i[24]&!i[23]&!i[22]
    &!i[21]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&i[30]&!i[29]
    &i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]&i[6]&!i[5]&i[4]&!i[3]
    &!i[2]&i[1]&i[0]) | (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]
    &!i[20]&!i[14]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&!i[26]
    &i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&i[12]&!i[6]&!i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]
    &!i[20]&i[13]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]
    &i[25]&i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[31]&!i[30]&!i[29]&i[28]&i[25]&i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&!i[29]&i[25]&i[14]&i[13]&!i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]
    &!i[27]&i[25]&i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]&i[25]&i[14]&!i[13]&!i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]&!i[14]&!i[6]
    &!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]&i[12]&!i[6]&!i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]&i[13]&!i[6]&!i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (i[15]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (i[16]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (i[17]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (i[18]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (i[19]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[14]&i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[14]&i[13]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[rs2] = (i[31]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[28]&i[27]&!i[26]&i[25]&!i[14]&!i[13]&!i[12]&!i[6]&!i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[28]&i[27]&!i[26]&i[25]&i[14]&i[13]&!i[6]&!i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[28]&i[27]&!i[26]&i[25]&i[14]&i[12]&!i[6]&!i[4]
    &!i[3]&i[2]&i[1]&i[0]);

assign out[rd] = (i[31]&i[29]&!i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]
    &!i[14]&!i[13]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&i[29]
    &!i[28]&!i[27]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&!i[14]&!i[13]
    &i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&i[30]&!i[29]&!i[28]
    &!i[27]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]&i[6]&!i[5]&i[4]&!i[3]&!i[2]
    &i[1]&i[0]) | (i[31]&i[30]&!i[29]&!i[28]&!i[27]&!i[26]&!i[24]&!i[23]
    &!i[22]&!i[21]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (i[14]&i[13]
    &i[12]&i[7]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[14]&i[13]
    &i[12]&i[8]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[14]&i[13]
    &i[12]&i[9]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[14]&i[13]
    &i[12]&i[10]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[14]&i[13]
    &i[12]&i[11]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]
    &i[29]&!i[28]&!i[27]&!i[25]&!i[14]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]
    &i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]&!i[27]&!i[26]&!i[14]&!i[13]
    &i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]
    &!i[27]&!i[26]&!i[14]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (
    i[31]&!i[30]&i[29]&!i[28]&!i[27]&!i[25]&!i[14]&!i[13]&i[6]&!i[5]&i[4]
    &!i[3]&!i[2]&i[1]&i[0]) | (i[15]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (i[16]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (i[17]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (i[18]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (i[19]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]);

assign out[vs1] = (!i[30]&!i[29]&i[28]&!i[27]&i[26]&i[25]&!i[14]&!i[13]&!i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[29]&!i[28]&i[26]&i[25]
    &!i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]
    &i[29]&!i[28]&i[27]&i[25]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[26]&!i[14]&!i[13]&i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]
    &!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]
    &!i[30]&!i[29]&i[25]&!i[14]&i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&i[30]&i[29]&!i[27]&i[25]&!i[14]&!i[13]&!i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&!i[28]
    &i[26]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[31]&!i[30]&!i[29]&i[28]&i[25]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&!i[27]&!i[26]&!i[14]
    &!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]
    &i[29]&!i[28]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]) | (i[31]&!i[30]&i[29]&!i[28]&!i[27]&i[25]&!i[14]&!i[13]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[30]&!i[29]&!i[27]&!i[26]
    &!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]
    &!i[30]&!i[29]&!i[26]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]&i[25]&!i[14]&!i[13]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vs2] = (!i[31]&!i[28]&!i[27]&!i[26]&!i[19]&!i[18]&!i[17]&!i[16]&!i[15]
    &!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[30]
    &!i[29]&i[28]&!i[27]&i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]&i[26]&i[25]&!i[14]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]
    &!i[27]&i[25]&!i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[31]&!i[30]&i[29]&!i[28]&i[27]&i[25]&!i[14]&i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[29]&!i[28]&i[27]&i[25]&!i[13]
    &!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]
    &!i[27]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]
    &i[29]&!i[28]&i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&!i[28]&i[27]&i[26]&!i[18]
    &!i[17]&!i[16]&!i[15]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[29]&!i[28]&i[27]&!i[26]&!i[19]&!i[18]&!i[17]
    &!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]
    &i[27]&i[26]&i[25]&i[14]&i[13]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[28]&i[27]&i[26]&i[25]&i[14]&i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[28]&i[27]&i[26]&i[25]&!i[14]&!i[13]&!i[12]&!i[6]&!i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (i[31]&!i[30]&!i[29]&i[25]&i[13]&!i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&!i[29]&i[28]&!i[27]&i[26]
    &i[25]&!i[14]&i[13]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]
    &i[30]&i[29]&i[28]&i[25]&!i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&i[25]&i[14]&!i[13]&!i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]&!i[27]
    &i[25]&!i[14]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]
    &i[30]&i[29]&!i[27]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&i[28]&i[25]&!i[13]&!i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[28]
    &!i[27]&!i[26]&i[25]&!i[14]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]) | (!i[31]&i[30]&i[29]&i[26]&i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]&!i[27]&i[25]
    &!i[13]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[30]&!i[29]&!i[27]
    &!i[26]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]
    &i[30]&i[29]&!i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]&i[25]&!i[13]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]&!i[13]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]
    &!i[28]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]
    &i[30]&i[29]&!i[28]&i[26]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]);

assign out[vs3] = (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&i[14]&i[13]
    &!i[6]&i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&!i[26]&i[25]&!i[24]
    &!i[23]&!i[22]&!i[21]&!i[20]&!i[14]&!i[13]&!i[12]&!i[6]&i[5]&!i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]
    &!i[21]&!i[20]&i[14]&i[12]&!i[6]&i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    i[31]&!i[30]&i[29]&!i[28]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[28]&i[27]&i[25]&i[14]&i[13]&!i[6]&i[5]&!i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]&!i[14]&!i[13]&!i[12]&!i[6]
    &i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]&i[14]&i[12]
    &!i[6]&i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vd] = (!i[30]&!i[29]&i[28]&!i[27]&i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&!i[27]&i[25]&!i[14]
    &i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[30]&i[29]
    &!i[28]&!i[27]&i[26]&i[25]&!i[14]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[30]&i[29]&!i[28]&i[27]&i[25]&!i[14]&i[13]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[29]&!i[28]
    &i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[31]&i[29]&!i[28]&i[27]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]&!i[13]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[28]
    &i[27]&i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&i[14]&!i[13]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&!i[26]&i[25]
    &!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&i[14]&i[13]&!i[6]&!i[5]&!i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]
    &!i[21]&!i[20]&i[14]&i[12]&!i[6]&!i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&!i[14]&!i[13]
    &!i[12]&!i[6]&!i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&!i[28]
    &i[27]&i[26]&!i[18]&!i[17]&!i[16]&!i[15]&!i[14]&!i[13]&i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[29]&!i[28]&i[27]&!i[26]
    &!i[19]&!i[18]&!i[17]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]
    &!i[20]&i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    i[31]&!i[30]&!i[29]&i[25]&i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&i[30]&i[29]&i[28]&i[25]&!i[14]&i[13]&i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&!i[29]&i[28]&!i[27]
    &i[26]&i[25]&!i[14]&i[13]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[28]&i[27]&i[25]&i[14]&i[13]&!i[6]&!i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[31]&i[30]&i[29]&i[25]&i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]&!i[27]&i[25]&!i[14]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]
    &!i[27]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[31]&!i[30]&!i[29]&i[28]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]&i[14]&i[12]&!i[6]&!i[5]&!i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&i[26]&i[14]&!i[13]&i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]&!i[14]
    &!i[13]&!i[12]&!i[6]&!i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]
    &i[29]&!i[28]&!i[27]&i[25]&!i[13]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]) | (!i[31]&!i[30]&!i[29]&!i[28]&!i[27]&!i[26]&i[25]&!i[14]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[30]&!i[29]&!i[27]
    &!i[26]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]
    &i[30]&i[29]&!i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]&!i[13]&i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]&i[25]&!i[13]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]
    &!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]
    &i[29]&!i[28]&i[26]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[imm12] = (!i[31]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[14]&i[13]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[14]&i[12]&!i[6]
    &!i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[simm] = (!i[30]&i[29]&!i[28]&!i[27]&i[26]&i[25]&!i[14]&i[13]&i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&!i[29]&i[28]&!i[27]
    &i[26]&i[25]&!i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[31]&!i[30]&!i[29]&!i[28]&!i[27]&!i[26]&i[25]&!i[14]&i[13]&i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&i[28]
    &i[25]&!i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    i[31]&!i[30]&i[29]&!i[28]&!i[27]&i[25]&!i[14]&i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&i[29]&!i[28]&i[27]&i[25]
    &!i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]
    &i[30]&i[29]&!i[27]&i[25]&!i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]);

assign out[vm ] = 1'b0;

assign out[vsetvl] = (i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[valu] = (!i[30]&i[29]&!i[28]&!i[27]&i[26]&i[25]&!i[14]&i[13]&i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[29]&!i[28]&i[26]&i[25]
    &!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[29]
    &!i[28]&i[27]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]) | (i[31]&!i[30]&!i[29]&i[28]&!i[27]&i[26]&i[25]&!i[14]&i[13]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]
    &!i[28]&!i[27]&i[25]&!i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&i[30]&i[29]&i[28]&i[25]&!i[14]&i[13]&i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[30]&!i[29]&i[28]&!i[27]&i[26]
    &i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]
    &!i[30]&!i[29]&!i[28]&!i[27]&!i[26]&i[25]&!i[14]&i[13]&i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&!i[27]&i[25]
    &!i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]
    &!i[30]&i[29]&!i[28]&i[27]&i[25]&!i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]&i[25]&!i[13]
    &!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]
    &i[28]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    i[31]&!i[30]&i[29]&!i[28]&!i[27]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&i[25]&i[14]&!i[13]&!i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&!i[27]
    &i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vmul] = (i[31]&!i[30]&!i[29]&i[28]&i[25]&i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]);

assign out[vdiv] = (i[31]&!i[30]&!i[29]&!i[28]&i[25]&i[13]&!i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]);

assign out[vrem] = (i[31]&!i[30]&!i[29]&!i[28]&i[27]&i[25]&i[13]&!i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vlsu] = (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&!i[14]
    &!i[13]&!i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&!i[26]
    &i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&i[14]&i[13]&!i[6]&!i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]
    &!i[21]&!i[20]&i[14]&i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[28]&i[27]&i[25]&!i[14]&!i[13]&!i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]
    &i[0]) | (!i[28]&i[27]&i[25]&i[14]&i[13]&!i[6]&!i[4]&!i[3]&i[2]&i[1]
    &i[0]) | (!i[28]&i[27]&i[25]&i[14]&i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]
    &i[0]);

assign out[vload] = (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&!i[14]
    &!i[13]&!i[12]&!i[6]&!i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]
    &!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&i[14]&i[13]&!i[6]
    &!i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&!i[26]&i[25]&!i[24]
    &!i[23]&!i[22]&!i[21]&!i[20]&i[14]&i[12]&!i[6]&!i[5]&!i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[28]&i[27]&i[25]&!i[14]&!i[13]&!i[12]&!i[6]&!i[5]
    &!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]&i[14]&i[13]&!i[6]
    &!i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]&i[14]&i[12]
    &!i[6]&!i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vstore] = (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&!i[14]
    &!i[13]&!i[12]&!i[6]&i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&!i[26]
    &i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&i[14]&i[13]&!i[6]&i[5]&!i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]
    &!i[21]&!i[20]&i[14]&i[12]&!i[6]&i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[28]&i[27]&i[25]&!i[14]&!i[13]&!i[12]&!i[6]&i[5]&!i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[28]&i[27]&i[25]&i[14]&i[13]&!i[6]&i[5]&!i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]&i[14]&i[12]&!i[6]&i[5]&!i[4]
    &!i[3]&i[2]&i[1]&i[0]);

assign out[vadd] = (!i[31]&!i[30]&!i[29]&!i[28]&!i[27]&!i[26]&i[25]&!i[14]&i[13]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]
    &!i[28]&!i[27]&!i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]);

assign out[vsub] = (!i[31]&i[30]&i[29]&!i[27]&i[25]&!i[14]&i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&i[28]&i[25]&!i[14]
    &i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]
    &!i[29]&i[27]&!i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&i[28]&i[25]&!i[13]&!i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&!i[28]&i[25]
    &!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]
    &i[29]&i[25]&i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[31]&i[30]&i[29]&!i[27]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]);

assign out[vand] = (!i[31]&!i[30]&i[29]&!i[28]&!i[27]&i[26]&i[25]&!i[14]&i[13]&i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&i[29]&!i[28]
    &!i[27]&i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]);

assign out[vor] = (!i[31]&!i[30]&i[29]&!i[28]&i[27]&!i[26]&i[25]&!i[14]&i[13]&i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&i[29]&!i[28]
    &i[27]&!i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]);

assign out[vxor] = (!i[31]&!i[30]&i[29]&!i[28]&i[27]&i[26]&i[25]&!i[14]&i[13]&i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&i[29]&!i[28]
    &i[27]&i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vsll] = (i[31]&!i[30]&!i[29]&i[28]&!i[27]&i[26]&i[25]&!i[14]&i[13]&i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&!i[29]&i[28]
    &!i[27]&i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]);

assign out[vsra] = (i[31]&!i[30]&i[29]&!i[28]&!i[27]&i[26]&i[25]&!i[14]&i[13]&i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]
    &!i[27]&i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]);

assign out[vsrl] = (i[31]&!i[30]&i[29]&!i[28]&!i[27]&!i[26]&i[25]&!i[14]&i[13]&i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]
    &!i[27]&!i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]);

assign out[vmslt] = (!i[31]&i[30]&i[29]&!i[28]&i[27]&i[25]&!i[13]&!i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vmseq] = (!i[31]&i[30]&i[29]&!i[28]&!i[27]&!i[26]&i[25]&!i[14]&i[13]&i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&!i[28]
    &!i[27]&!i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]);

assign out[vmsne] = (!i[31]&i[30]&i[29]&!i[28]&!i[27]&i[26]&i[25]&!i[14]&i[13]&i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&!i[28]
    &!i[27]&i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]);

assign out[vmsle] = (!i[31]&i[30]&i[29]&i[28]&!i[27]&i[25]&!i[14]&i[13]&i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&i[28]&!i[27]
    &i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vmsgt] = (!i[31]&i[30]&i[29]&i[28]&i[27]&i[25]&i[14]&!i[13]&!i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&i[28]&i[27]
    &i[25]&!i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[unsign] = (!i[31]&i[30]&i[29]&i[27]&!i[26]&i[25]&i[14]&!i[13]&!i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&!i[29]&!i[28]&i[27]
    &!i[26]&!i[19]&!i[18]&!i[17]&!i[15]&!i[14]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&i[30]&!i[29]&!i[27]&!i[25]&!i[24]
    &!i[23]&!i[22]&!i[21]&i[20]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (
    i[31]&i[30]&!i[29]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]&i[20]
    &i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&i[28]
    &!i[26]&i[25]&!i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[31]&i[30]&i[29]&!i[28]&i[27]&!i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&!i[29]&!i[26]&i[25]&i[13]
    &!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]
    &i[28]&!i[27]&!i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&i[28]&!i[26]&i[25]&!i[13]&!i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[sign] = (!i[31]&i[30]&i[29]&i[27]&i[26]&i[25]&i[14]&!i[13]&!i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&!i[29]&!i[28]&i[27]
    &!i[26]&!i[19]&!i[18]&!i[17]&i[15]&!i[14]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&i[30]&!i[29]&!i[27]&!i[25]&!i[24]
    &!i[23]&!i[22]&!i[21]&!i[20]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (
    i[31]&i[30]&!i[29]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]
    &i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&i[28]
    &i[26]&i[25]&!i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[31]&i[30]&i[29]&!i[28]&i[27]&i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&!i[29]&i[26]&i[25]&i[13]
    &!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]
    &i[28]&!i[27]&i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&i[28]&i[26]&i[25]&!i[13]&!i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[by] = (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&!i[14]&!i[13]
    &!i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]&!i[14]
    &!i[13]&!i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[half] = (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&i[14]
    &!i[13]&i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]
    &i[14]&!i[13]&i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[word] = (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&i[14]
    &i[13]&!i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]
    &i[14]&i[13]&!i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[element] = (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&i[14]
    &i[13]&i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]
    &i[14]&i[13]&i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[csr_read] = (!i[19]&!i[18]&!i[17]&!i[16]&!i[15]&i[14]&i[13]&i[12]&!i[11]
    &!i[10]&!i[9]&!i[8]&!i[7]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[csr_write_1] = (i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[csr_write_2] = (i[14]&i[13]&i[12]&i[7]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]) | (i[14]&i[13]&i[12]&i[8]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    i[14]&i[13]&i[12]&i[9]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    i[14]&i[13]&i[12]&i[10]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    i[14]&i[13]&i[12]&i[11]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    i[15]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    i[16]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    i[17]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    i[18]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    i[19]&i[14]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[rs1_sign] = (i[31]&!i[30]&!i[29]&i[28]&i[27]&i[26]&i[25]&i[14]&i[13]&!i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[rs2_sign ] = 1'b0;

assign out[vs1_sign] = (i[31]&!i[30]&!i[29]&i[28]&i[27]&i[26]&i[25]&!i[14]&i[13]
    &!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vs2_sign] = (i[31]&!i[30]&!i[29]&i[28]&i[27]&i[25]&i[13]&!i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[low] = (i[31]&!i[30]&!i[29]&i[28]&!i[27]&i[26]&i[25]&i[13]&!i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[unit_st] = (!i[28]&!i[27]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]
    &!i[14]&!i[13]&!i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]
    &!i[27]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&i[14]&i[13]
    &!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&!i[27]&!i[26]&i[25]
    &!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&i[14]&i[12]&!i[6]&!i[4]&!i[3]
    &i[2]&i[1]&i[0]);

assign out[stride] = (!i[28]&i[27]&!i[26]&i[25]&!i[14]&!i[13]&!i[12]&!i[6]&!i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[28]&i[27]&!i[26]&i[25]&i[14]&i[13]&!i[6]&!i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (!i[28]&i[27]&!i[26]&i[25]&i[14]&i[12]&!i[6]
    &!i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[indexed] = (!i[28]&i[27]&i[26]&i[25]&!i[14]&!i[13]&!i[12]&!i[6]&!i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[26]&i[25]&i[14]&i[13]&!i[6]&!i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[26]&i[25]&i[14]&i[12]&!i[6]
    &!i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[zero_extend] = (i[31]&!i[30]&!i[29]&i[28]&!i[27]&i[26]&i[25]&!i[14]&i[13]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]
    &!i[28]&!i[27]&!i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]&!i[27]&i[25]&!i[14]&i[13]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[sign_extend] = (i[31]&!i[30]&!i[29]&i[28]&!i[27]&i[26]&i[25]&!i[13]&!i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&!i[26]&i[25]&!i[24]
    &!i[23]&!i[22]&!i[21]&!i[20]&i[14]&i[13]&!i[6]&!i[5]&!i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]
    &!i[14]&!i[13]&!i[12]&!i[6]&!i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&i[14]&i[12]
    &!i[6]&!i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]
    &!i[27]&i[26]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]) | (!i[28]&i[27]&i[25]&i[14]&i[13]&!i[6]&!i[5]&!i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[28]&i[27]&i[25]&!i[14]&!i[13]&!i[12]&!i[6]&!i[5]
    &!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]&i[14]&i[12]&!i[6]
    &!i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[i0_only] = (i[31]&!i[30]&!i[29]&!i[28]&i[25]&i[13]&!i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]);

assign out[vmin] = (!i[31]&!i[30]&!i[29]&i[28]&!i[27]&i[25]&!i[13]&!i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vmax] = (!i[31]&!i[30]&!i[29]&i[28]&i[27]&i[25]&!i[13]&!i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[fs1] = (i[31]&i[29]&!i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]
    &!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&i[29]&!i[28]
    &!i[27]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&!i[14]&!i[13]&i[6]
    &!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[26]&i[14]
    &!i[13]&i[12]&i[6]&!i[5]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]
    &!i[27]&i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[30]&i[29]&!i[28]&!i[27]&i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[28]&i[27]&i[26]&i[25]&!i[24]&!i[23]
    &!i[22]&!i[21]&!i[20]&i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]
    &!i[20]&i[14]&!i[13]&i[12]&i[6]&!i[5]&!i[3]&i[2]&i[1]&i[0]) | (i[31]
    &i[30]&!i[29]&!i[28]&!i[27]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]&i[6]
    &!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&i[30]&!i[29]&!i[28]&!i[27]
    &!i[26]&!i[24]&!i[23]&!i[22]&!i[21]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[31]&i[30]&i[29]&i[26]&i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]&!i[25]&!i[14]&!i[12]
    &i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]
    &!i[26]&!i[14]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]
    &!i[30]&!i[29]&!i[26]&i[14]&!i[13]&i[12]&i[6]&!i[5]&!i[3]&i[1]&i[0]) | (
    !i[30]&!i[29]&!i[27]&!i[26]&i[14]&!i[13]&i[12]&i[6]&!i[5]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[30]&!i[28]&!i[25]&!i[14]&!i[13]&i[6]&!i[5]
    &!i[3]&!i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]&i[14]&!i[13]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[28]
    &!i[26]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[30]
    &i[29]&!i[28]&!i[27]&!i[25]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]
    &i[0]) | (!i[30]&i[29]&!i[28]&!i[27]&!i[26]&!i[14]&!i[13]&i[6]&!i[5]
    &!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[29]&i[28]&i[27]&!i[25]&i[6]&!i[5]
    &!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[29]&i[28]&i[27]&!i[26]&i[6]&!i[5]
    &!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[25]&i[6]&!i[5]
    &!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]&i[6]&!i[5]
    &!i[3]&!i[2]&i[1]&i[0]) | (!i[25]&i[6]&!i[5]&!i[4]&i[1]&i[0]) | (
    !i[26]&i[6]&!i[5]&!i[4]&i[1]&i[0]);

assign out[fs2] = (!i[30]&i[29]&!i[28]&!i[27]&!i[25]&!i[14]&!i[12]&i[6]&!i[5]&!i[3]
    &!i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]&!i[26]&!i[14]&!i[12]
    &i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]
    &!i[25]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[30]
    &i[29]&!i[28]&!i[27]&!i[26]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]
    &i[0]) | (!i[31]&!i[30]&!i[28]&!i[25]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]
    &!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[28]&!i[26]&!i[14]&!i[13]&i[6]
    &!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[14]&i[13]&!i[6]&i[5]&!i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[14]&i[12]&!i[6]&i[5]&!i[4]&!i[3]&i[2]&i[1]
    &i[0]) | (!i[31]&!i[30]&!i[29]&!i[25]&i[6]&!i[5]&!i[3]&!i[2]&i[1]
    &i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]&i[6]&!i[5]&!i[3]&!i[2]&i[1]
    &i[0]) | (!i[25]&i[6]&!i[5]&!i[4]&i[1]&i[0]) | (!i[26]&i[6]&!i[5]
    &!i[4]&i[1]&i[0]);

assign out[fs3] = (!i[25]&i[6]&!i[5]&!i[4]&i[1]&i[0]) | (!i[26]&i[6]&!i[5]&!i[4]&i[1]
    &i[0]);

assign out[fd] = (!i[31]&i[30]&!i[29]&!i[28]&!i[27]&!i[26]&!i[19]&!i[18]&!i[17]&!i[16]
    &!i[15]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&!i[3]&i[2]&i[1]&i[0]) | (
    i[31]&i[30]&i[28]&!i[27]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]
    &!i[14]&!i[13]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]
    &i[30]&i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&!i[14]
    &!i[13]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&i[30]&!i[29]
    &i[28]&!i[27]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]&i[6]&!i[5]&!i[3]
    &!i[2]&i[1]&i[0]) | (i[31]&i[30]&!i[29]&i[28]&!i[27]&!i[26]&!i[24]
    &!i[23]&!i[22]&!i[21]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]
    &!i[30]&!i[28]&!i[25]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[31]&!i[30]&!i[28]&!i[26]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]
    &i[0]) | (!i[31]&!i[30]&!i[28]&!i[27]&!i[25]&!i[14]&!i[12]&i[6]&!i[5]
    &!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[28]&!i[27]&!i[26]&!i[14]
    &!i[12]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[14]&i[13]&!i[6]&!i[5]
    &!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[29]&i[28]&i[27]&!i[25]&i[6]
    &!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[29]&i[28]&i[27]&!i[26]
    &i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[14]&i[12]&!i[6]&!i[5]&!i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[25]&i[6]&!i[5]&!i[3]
    &!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]&i[6]&!i[5]&!i[3]
    &!i[2]&i[1]&i[0]) | (!i[25]&i[6]&!i[5]&!i[4]&i[1]&i[0]) | (!i[26]
    &i[6]&!i[5]&!i[4]&i[1]&i[0]);

assign out[vfadd] = (!i[31]&!i[30]&!i[29]&!i[28]&!i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfsub] = (!i[31]&!i[30]&!i[29]&!i[28]&i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfmin] = (!i[31]&!i[30]&!i[29]&i[28]&!i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfmax] = (!i[31]&!i[30]&!i[29]&i[28]&i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfmv] = (!i[31]&i[30]&!i[29]&i[28]&i[27]&i[26]&i[25]&!i[24]&!i[23]&!i[22]
    &!i[21]&!i[20]&i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]);

assign out[vfmvs] = (!i[31]&i[30]&!i[29]&!i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]
    &!i[21]&!i[20]&i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]);

assign out[vfmvf] = (!i[31]&i[30]&!i[29]&!i[28]&!i[27]&!i[26]&!i[19]&!i[18]&!i[17]
    &!i[16]&!i[15]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]);

assign out[vmfeq] = (!i[31]&i[30]&i[29]&!i[28]&!i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vmfle] = (!i[31]&i[30]&i[29]&!i[28]&!i[27]&i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vmflt] = (!i[31]&i[30]&i[29]&!i[28]&i[27]&i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vmfne] = (!i[31]&i[30]&i[29]&i[28]&!i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vmfgt] = (!i[31]&i[30]&i[29]&i[28]&!i[27]&i[26]&i[14]&!i[13]&i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vmfge] = (!i[31]&i[30]&i[29]&i[28]&i[27]&i[26]&i[14]&!i[13]&i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfdiv] = (i[31]&!i[30]&!i[29]&!i[28]&!i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfmul] = (i[31]&!i[30]&!i[29]&i[28]&!i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfmadd] = (i[31]&!i[30]&i[29]&!i[28]&!i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfmsub] = (i[31]&!i[30]&i[29]&!i[28]&i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfnmadd] = (i[31]&!i[30]&i[29]&!i[28]&!i[27]&i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfnmsub] = (i[31]&!i[30]&i[29]&!i[28]&i[27]&i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfsqrt] = (!i[31]&i[30]&!i[29]&!i[28]&i[27]&i[26]&!i[19]&!i[18]&!i[17]
    &!i[16]&!i[15]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]);

assign out[vfcvt_x_f] = (!i[31]&i[30]&!i[29]&!i[28]&i[27]&!i[26]&!i[19]&!i[18]&!i[17]
    &!i[16]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfcvt_f_x] = (!i[31]&i[30]&!i[29]&!i[28]&i[27]&!i[26]&!i[19]&!i[18]&!i[17]
    &i[16]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfsgnj] = (!i[31]&!i[30]&i[29]&!i[28]&!i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfsgnjn] = (!i[31]&!i[30]&i[29]&!i[28]&!i[27]&i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfsgnjx] = (!i[31]&!i[30]&i[29]&!i[28]&i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[vfclass] = (!i[31]&i[30]&!i[29]&!i[28]&i[27]&i[26]&i[19]&!i[18]&!i[17]
    &!i[16]&!i[15]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]);

assign out[vfpu] = (!i[31]&!i[28]&!i[27]&!i[26]&!i[19]&!i[18]&!i[17]&!i[16]&!i[15]
    &!i[14]&!i[13]&i[12]&i[6]&!i[5]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&i[29]
    &!i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&!i[14]&!i[13]
    &i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&i[29]&!i[28]&!i[27]&!i[25]
    &!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]
    &!i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]&!i[26]&!i[14]&!i[13]
    &i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[26]
    &!i[13]&i[12]&i[6]&!i[5]&!i[3]&i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]
    &!i[27]&!i[25]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[30]&i[29]&!i[28]&!i[27]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&i[30]&i[28]&i[27]&i[26]&i[25]&!i[24]&!i[23]
    &!i[22]&!i[21]&!i[20]&i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (i[31]&i[30]&!i[27]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]
    &!i[20]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    i[31]&i[30]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&!i[14]
    &!i[13]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&i[30]
    &!i[28]&i[27]&i[26]&!i[18]&!i[17]&!i[16]&!i[15]&!i[14]&!i[13]&i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[29]&!i[28]&i[27]
    &!i[26]&!i[19]&!i[18]&!i[17]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[31]&!i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]
    &!i[21]&!i[20]&i[14]&!i[13]&i[12]&i[6]&!i[5]&!i[3]&i[2]&i[1]&i[0]) | (
    i[31]&i[30]&!i[29]&!i[27]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]&i[6]
    &!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&i[30]&!i[29]&!i[27]&!i[26]
    &!i[24]&!i[23]&!i[22]&!i[21]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[30]&i[29]&!i[28]&!i[27]&!i[25]&!i[14]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]
    &i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]&!i[26]&!i[14]&!i[12]&i[6]
    &!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&i[26]&i[14]&!i[13]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[28]
    &!i[25]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]
    &!i[30]&!i[28]&!i[26]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    i[31]&!i[30]&i[29]&!i[28]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &!i[3]&i[1]&i[0]) | (!i[30]&!i[29]&!i[27]&!i[26]&!i[13]&i[12]&i[6]
    &!i[5]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&!i[27]&!i[26]
    &!i[13]&i[12]&i[6]&!i[5]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]
    &!i[28]&i[26]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[31]&!i[29]&i[28]&i[27]&!i[25]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[31]&!i[29]&i[28]&i[27]&!i[26]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[31]&!i[30]&!i[29]&!i[25]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[31]&!i[30]&!i[29]&!i[26]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[25]&i[6]&!i[5]&!i[4]&i[1]&i[0]) | (!i[26]&i[6]&!i[5]&!i[4]&i[1]
    &i[0]);

assign out[fadd] = (!i[31]&!i[30]&!i[29]&!i[28]&!i[27]&!i[25]&i[6]&!i[5]&i[4]&!i[3]
    &!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[28]&!i[27]&!i[26]&i[6]
    &!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]);

assign out[fsub] = (!i[31]&!i[30]&!i[29]&!i[28]&i[27]&!i[25]&i[6]&!i[5]&i[4]&!i[3]
    &!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[28]&i[27]&!i[26]&i[6]
    &!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]);

assign out[fmul] = (!i[31]&!i[30]&!i[29]&i[28]&!i[27]&!i[25]&i[6]&!i[5]&i[4]&!i[3]
    &!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&i[28]&!i[27]&!i[26]&i[6]
    &!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]);

assign out[fdiv] = (!i[31]&!i[30]&!i[29]&i[28]&i[27]&!i[25]&i[6]&!i[5]&i[4]&!i[3]
    &!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&i[28]&i[27]&!i[26]&i[6]
    &!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]);

assign out[fsqrt] = (!i[31]&i[30]&!i[29]&i[28]&i[27]&!i[25]&i[6]&!i[5]&i[4]&!i[3]
    &!i[2]&i[1]&i[0]) | (!i[31]&i[30]&!i[29]&i[28]&i[27]&!i[26]&i[6]&!i[5]
    &i[4]&!i[3]&!i[2]&i[1]&i[0]);

assign out[fmin] = (!i[31]&!i[30]&i[29]&!i[28]&i[27]&!i[25]&!i[14]&!i[13]&!i[12]&i[6]
    &!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&i[29]&!i[28]
    &i[27]&!i[26]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]
    &i[0]);

assign out[fmax] = (!i[31]&!i[30]&i[29]&!i[28]&i[27]&!i[25]&!i[14]&!i[13]&i[12]&i[6]
    &!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&i[29]&!i[28]
    &i[27]&!i[26]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]
    &i[0]);

assign out[fmvx] = (i[31]&i[30]&i[29]&i[28]&!i[27]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]
    &!i[20]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (
    i[31]&i[30]&i[29]&i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]
    &!i[20]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]);

assign out[fmvf] = (i[31]&i[30]&i[29]&!i[28]&!i[27]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]
    &!i[20]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (
    i[31]&i[30]&i[29]&!i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]
    &!i[20]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]);

assign out[feq] = (i[31]&!i[30]&i[29]&!i[28]&!i[27]&!i[25]&!i[14]&i[13]&!i[12]&i[6]
    &!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]&!i[27]
    &!i[26]&!i[14]&i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]);

assign out[flt] = (i[31]&!i[30]&i[29]&!i[28]&!i[27]&!i[25]&!i[14]&!i[13]&i[12]&i[6]
    &!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]&!i[27]
    &!i[26]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]);

assign out[fle] = (i[31]&!i[30]&i[29]&!i[28]&!i[27]&!i[25]&!i[14]&!i[13]&!i[12]&i[6]
    &!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]&!i[27]
    &!i[26]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]);

assign out[fmadd] = (!i[25]&i[6]&!i[5]&!i[4]&!i[3]&!i[2]&i[1]&i[0]) | (!i[26]&i[6]
    &!i[5]&!i[4]&!i[3]&!i[2]&i[1]&i[0]);

assign out[fmsub] = (!i[25]&i[6]&!i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[26]&i[6]
    &!i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[fnmsub] = (!i[25]&i[6]&!i[5]&!i[4]&i[3]&!i[2]&i[1]&i[0]) | (!i[26]&i[6]
    &!i[5]&!i[4]&i[3]&!i[2]&i[1]&i[0]);

assign out[fnmadd] = (!i[25]&i[6]&!i[5]&!i[4]&i[3]&i[2]&i[1]&i[0]) | (!i[26]&i[6]
    &!i[5]&!i[4]&i[3]&i[2]&i[1]&i[0]);

assign out[fsgnj] = (!i[31]&!i[30]&i[29]&!i[28]&!i[27]&!i[25]&!i[14]&!i[13]&!i[12]
    &i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&i[29]&!i[28]
    &!i[27]&!i[26]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]
    &i[0]);

assign out[fsgnjn] = (!i[31]&!i[30]&i[29]&!i[28]&!i[27]&!i[25]&!i[14]&!i[13]&i[12]
    &i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&i[29]&!i[28]
    &!i[27]&!i[26]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]
    &i[0]);

assign out[fsgnjx] = (!i[31]&!i[30]&i[29]&!i[28]&!i[27]&!i[25]&!i[14]&i[13]&!i[12]
    &i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&i[29]&!i[28]
    &!i[27]&!i[26]&!i[14]&i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]
    &i[0]);

assign out[fcvt_w_p] = (i[31]&i[30]&!i[29]&!i[28]&!i[27]&!i[25]&!i[24]&!i[23]&!i[22]
    &!i[21]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&i[30]&!i[29]
    &!i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]&i[6]&!i[5]&i[4]
    &!i[3]&!i[2]&i[1]&i[0]);

assign out[fcvt_p_w] = (i[31]&i[30]&!i[29]&i[28]&!i[27]&!i[25]&!i[24]&!i[23]&!i[22]
    &!i[21]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&i[30]&!i[29]
    &i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]&i[6]&!i[5]&i[4]&!i[3]
    &!i[2]&i[1]&i[0]);

assign out[fclass] = (i[31]&i[30]&i[29]&!i[28]&!i[27]&!i[25]&!i[24]&!i[23]&!i[22]
    &!i[21]&!i[20]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]
    &i[0]) | (i[31]&i[30]&i[29]&!i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]
    &!i[21]&!i[20]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&!i[2]&i[1]
    &i[0]);

assign out[flsu] = (!i[14]&i[13]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[14]&i[12]
    &!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[fload] = (!i[14]&i[13]&!i[6]&!i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[14]
    &i[12]&!i[6]&!i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[fstore] = (!i[14]&i[13]&!i[6]&i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[14]
    &i[12]&!i[6]&i[5]&!i[4]&!i[3]&i[2]&i[1]&i[0]);

assign out[single_p] = (i[31]&i[29]&!i[28]&!i[27]&!i[26]&!i[25]&!i[24]&!i[23]&!i[22]
    &!i[21]&!i[20]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    i[31]&i[30]&!i[27]&!i[26]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]
    &!i[14]&!i[13]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]
    &i[30]&!i[29]&!i[27]&!i[26]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]&i[6]
    &!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[28]&!i[26]&!i[25]
    &!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[14]&i[13]
    &!i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]
    &!i[27]&!i[26]&!i[25]&!i[14]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[30]&i[29]&!i[28]&!i[27]&!i[26]&!i[25]&!i[14]&!i[13]&i[6]&!i[5]
    &!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[29]&i[28]&i[27]&!i[26]&!i[25]
    &i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]
    &!i[25]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[26]&!i[25]&i[6]&!i[5]
    &!i[4]&i[1]&i[0]);

assign out[double_p] = (i[31]&i[29]&!i[28]&!i[27]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]
    &!i[21]&!i[20]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    i[31]&i[30]&!i[27]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]
    &!i[14]&!i[13]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]
    &i[30]&!i[29]&!i[27]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&i[6]
    &!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[14]&i[13]&i[12]&!i[6]&!i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[28]&!i[26]&i[25]&!i[14]&!i[13]
    &i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]
    &!i[26]&i[25]&!i[14]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[30]&i[29]&!i[28]&!i[27]&!i[26]&i[25]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]
    &!i[2]&i[1]&i[0]) | (!i[31]&!i[29]&i[28]&i[27]&!i[26]&i[25]&i[6]&!i[5]
    &!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]&i[25]&i[6]
    &!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[26]&i[25]&i[6]&!i[5]&!i[4]&i[1]
    &i[0]);

assign out[half_p] = (i[31]&i[29]&!i[28]&!i[27]&i[26]&!i[25]&!i[24]&!i[23]&!i[22]
    &!i[21]&!i[20]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    i[31]&i[30]&!i[27]&i[26]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]
    &!i[14]&!i[13]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]
    &i[30]&!i[29]&!i[27]&i[26]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]&i[6]
    &!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[28]&i[26]&!i[25]
    &!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[30]&i[29]
    &!i[28]&!i[27]&i[26]&!i[25]&!i[14]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]&i[1]
    &i[0]) | (!i[14]&!i[13]&i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[30]&i[29]&!i[28]&!i[27]&i[26]&!i[25]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]
    &!i[2]&i[1]&i[0]) | (!i[31]&!i[29]&i[28]&i[27]&i[26]&!i[25]&i[6]&!i[5]
    &!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&i[26]&!i[25]&i[6]
    &!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (i[26]&!i[25]&i[6]&!i[5]&!i[4]&i[1]
    &i[0]);

assign out[scalar_fpu] = (i[31]&i[29]&!i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]
    &!i[20]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]
    &i[29]&!i[28]&!i[27]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&!i[14]
    &!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&i[30]&!i[27]&!i[25]
    &!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]
    &!i[3]&!i[2]&i[1]&i[0]) | (i[31]&i[30]&!i[27]&!i[26]&!i[24]&!i[23]
    &!i[22]&!i[21]&!i[20]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]
    &i[1]&i[0]) | (i[31]&i[30]&!i[29]&!i[27]&!i[25]&!i[24]&!i[23]&!i[22]
    &!i[21]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (i[31]&i[30]&!i[29]&!i[27]
    &!i[26]&!i[24]&!i[23]&!i[22]&!i[21]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[31]&!i[30]&!i[28]&!i[25]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]
    &i[0]) | (!i[31]&!i[30]&!i[28]&!i[26]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]
    &!i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]&!i[25]&!i[14]&!i[12]
    &i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]
    &!i[26]&!i[14]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[30]
    &i[29]&!i[28]&!i[27]&!i[25]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]
    &i[0]) | (!i[30]&i[29]&!i[28]&!i[27]&!i[26]&!i[14]&!i[13]&i[6]&!i[5]
    &!i[3]&!i[2]&i[1]&i[0]) | (!i[14]&i[13]&!i[6]&!i[4]&!i[3]&i[2]&i[1]
    &i[0]) | (!i[14]&i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]
    &!i[29]&i[28]&i[27]&!i[25]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[31]&!i[29]&i[28]&i[27]&!i[26]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[31]&!i[30]&!i[29]&!i[25]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[31]&!i[30]&!i[29]&!i[26]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[25]&i[6]&!i[5]&!i[4]&i[1]&i[0]) | (!i[26]&i[6]&!i[5]&!i[4]&i[1]
    &i[0]);

assign out[vector_fpu] = (!i[31]&!i[28]&!i[27]&!i[26]&!i[19]&!i[18]&!i[17]&!i[16]
    &!i[15]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[30]&i[29]&!i[28]&!i[27]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[26]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[28]&i[27]&i[26]&i[25]
    &!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&i[14]&!i[13]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&!i[28]&i[27]&i[26]&!i[18]
    &!i[17]&!i[16]&!i[15]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]
    &!i[20]&i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[31]&!i[29]&!i[28]&i[27]&!i[26]&!i[19]&!i[18]&!i[17]&!i[14]&!i[13]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]
    &i[26]&i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[30]&!i[29]&!i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (i[31]&!i[30]&i[29]&!i[28]&!i[13]&i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]&!i[13]&i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&!i[27]
    &!i[26]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]
    &i[30]&i[29]&!i[28]&i[26]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]);

assign out[legal] = (i[31]&i[29]&!i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]
    &!i[20]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]
    &!i[28]&!i[27]&!i[26]&!i[19]&!i[18]&!i[17]&!i[16]&!i[15]&!i[14]&!i[13]
    &i[12]&i[6]&!i[5]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&i[29]&!i[28]&!i[27]
    &!i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&!i[14]&!i[13]&i[6]&!i[5]
    &!i[3]&!i[2]&i[1]&i[0]) | (!i[30]&!i[29]&i[28]&!i[27]&i[26]&i[25]
    &!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]
    &i[29]&i[25]&i[14]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    i[31]&!i[30]&i[29]&!i[28]&!i[27]&i[25]&i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&i[26]&i[14]&i[12]&i[6]&!i[5]
    &i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]&!i[25]
    &!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&!i[30]
    &!i[28]&!i[26]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (
    !i[31]&!i[30]&i[29]&!i[28]&i[27]&i[25]&i[13]&i[12]&i[6]&!i[5]&i[4]
    &!i[3]&i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]&i[26]&i[25]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&i[29]
    &!i[28]&!i[27]&i[25]&!i[13]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[31]&i[30]&i[29]&!i[27]&i[25]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]&!i[26]&!i[14]&!i[13]
    &i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]
    &i[26]&i[25]&!i[13]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[30]
    &i[29]&!i[28]&!i[26]&!i[13]&i[12]&i[6]&!i[5]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[31]&i[29]&!i[28]&i[27]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[31]&i[30]&i[29]&!i[28]&i[26]&!i[13]&i[12]&i[6]
    &!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]&!i[13]
    &i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[14]&i[13]&i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&i[30]&!i[27]&!i[25]
    &!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]
    &!i[3]&!i[2]&i[1]&i[0]) | (i[31]&i[30]&!i[27]&!i[26]&!i[24]&!i[23]
    &!i[22]&!i[21]&!i[20]&!i[14]&!i[13]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]
    &i[1]&i[0]) | (!i[31]&i[30]&i[28]&i[27]&i[26]&i[25]&!i[24]&!i[23]
    &!i[22]&!i[21]&!i[20]&i[14]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]) | (!i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]
    &i[13]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[28]&!i[26]&i[25]&!i[24]
    &!i[23]&!i[22]&!i[21]&!i[20]&!i[14]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[28]&!i[26]&i[25]&!i[24]&!i[23]&!i[22]&!i[21]&!i[20]&i[12]&!i[6]
    &!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&i[30]&!i[28]&i[27]&i[26]&!i[18]
    &!i[17]&!i[16]&!i[15]&!i[14]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[29]&!i[28]&i[27]&!i[26]&!i[19]&!i[18]&!i[17]
    &!i[14]&!i[13]&i[12]&i[6]&!i[5]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&i[30]
    &!i[29]&!i[27]&!i[25]&!i[24]&!i[23]&!i[22]&!i[21]&i[6]&!i[5]&!i[3]
    &!i[2]&i[1]&i[0]) | (!i[31]&!i[28]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]
    &!i[21]&!i[20]&i[14]&i[12]&i[6]&!i[5]&!i[3]&i[2]&i[1]&i[0]) | (i[31]
    &i[30]&!i[29]&!i[27]&!i[26]&!i[24]&!i[23]&!i[22]&!i[21]&i[6]&!i[5]
    &!i[3]&!i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]&!i[25]&!i[14]
    &!i[12]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[28]&i[27]&i[25]&i[13]
    &!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]&!i[30]&!i[29]&i[25]&i[13]
    &!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[28]
    &!i[25]&!i[14]&!i[13]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]
    &i[30]&i[29]&i[28]&i[25]&i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]
    &i[0]) | (!i[28]&i[27]&i[25]&!i[14]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[28]&i[27]&i[25]&i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (i[31]
    &!i[30]&!i[29]&i[28]&!i[27]&i[26]&i[25]&i[13]&i[6]&!i[5]&i[4]&!i[3]
    &i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&i[28]&i[25]&!i[13]&!i[12]
    &i[6]&!i[5]&i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[30]&i[29]&!i[28]&!i[27]
    &!i[26]&!i[14]&!i[12]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]
    &i[30]&i[29]&!i[27]&i[25]&!i[13]&!i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]&i[25]&!i[13]&i[6]&!i[5]
    &!i[3]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[28]&!i[27]&!i[26]&i[25]
    &i[12]&i[6]&!i[5]&!i[3]&i[1]&i[0]) | (!i[30]&!i[29]&!i[27]&!i[26]
    &!i[13]&i[12]&i[6]&!i[5]&!i[3]&i[2]&i[1]&i[0]) | (!i[31]&!i[30]&!i[29]
    &!i[26]&!i[13]&i[12]&i[6]&!i[5]&!i[3]&i[1]&i[0]) | (!i[31]&!i[29]
    &i[28]&i[27]&!i[25]&i[6]&!i[5]&!i[3]&!i[2]&i[1]&i[0]) | (!i[31]&i[30]
    &i[29]&!i[27]&!i[26]&!i[13]&i[12]&i[6]&!i[5]&!i[3]&i[2]&i[1]&i[0]) | (
    i[31]&!i[30]&i[29]&!i[28]&!i[13]&i[12]&i[6]&!i[5]&i[4]&!i[3]&i[2]
    &i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[25]&i[6]&!i[5]&!i[3]&!i[2]
    &i[1]&i[0]) | (!i[31]&!i[29]&i[28]&i[27]&!i[26]&i[6]&!i[5]&!i[3]&!i[2]
    &i[1]&i[0]) | (!i[31]&!i[30]&!i[29]&!i[26]&i[6]&!i[5]&!i[3]&!i[2]
    &i[1]&i[0]) | (!i[14]&i[13]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (
    !i[14]&i[12]&!i[6]&!i[4]&!i[3]&i[2]&i[1]&i[0]) | (!i[25]&i[6]&!i[5]
    &!i[4]&i[1]&i[0]) | (!i[26]&i[6]&!i[5]&!i[4]&i[1]&i[0]);





endmodule
