module FPU_move(rst_l,opcode,Move_Input_IEEE,Move_Output_IEEE);
  //Standard Defination For Parameterization
  
  parameter Std = 31; // Means IEEE754 Std 32 Bit Single Precision -1 for bits
  
  input [Std : 0] Move_Input_IEEE; // Input of IEEE754 32 Move Instruction 
  input [1:0] opcode; // opcode for selection
  input rst_l; // clock & reset for Synchronizations
  output [Std : 0] Move_Output_IEEE; // Output of IEEE754 32 Move Instruction 
  
  wire [Std : 0] Move_Output_IEEE; // Define reg becuase it is Output of IEEE754 32 Move Instruction 
   
  // New logic will  be
  assign Move_Output_IEEE = (rst_l == 1'b0) ? 32'h00000000 :  (opcode[0] == 1'b1) ? Move_Input_IEEE : (opcode[1] == 1'b1) ? Move_Input_IEEE : 32'h00000000;
  
endmodule
